----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    14:54:38 05/21/2015 
-- Design Name: 
-- Module Name:    ItoA - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity ItoA is
    Port ( I : in  STD_LOGIC_VECTOR (7 downto 0);
           A : out  STD_LOGIC_VECTOR (31 downto 0);
			  l : out integer);
end ItoA;

architecture Behavioral of ItoA is

begin


ITOA: process(I)
begin

		case I is 
			 when X"00" =>  A <= X"20202030"; -- 000
							 l <= 2;
			 when X"01" =>  A <= X"20202031"; -- 001
							 l <= 2;
			 when X"02" =>  A <= X"20202032"; -- 002
							 l <= 2;
			 when X"03" =>  A <= X"20202033"; -- 003
							 l <= 2;
			 when X"04" =>  A <= X"20202034"; -- 004
							 l <= 2;
			 when X"05" =>  A <= X"20202035"; -- 005
							 l <= 2;
			 when X"06" =>  A <= X"20202036"; -- 006
							 l <= 2;
			 when X"07" =>  A <= X"20202037"; -- 007
							 l <= 2;
			 when X"08" =>  A <= X"20202038"; -- 008
							 l <= 2;
			 when X"09" =>  A <= X"20202039"; -- 009
							 l <= 2;
			 when X"0a" =>  A <= X"20203130"; -- 010
							 l <= 3;
			 when X"0b" =>  A <= X"20203131"; -- 011
							 l <= 3;
			 when X"0c" =>  A <= X"20203132"; -- 012
							 l <= 3;
			 when X"0d" =>  A <= X"20203133"; -- 013
							 l <= 3;
			 when X"0e" =>  A <= X"20203134"; -- 014
							 l <= 3;
			 when X"0f" =>  A <= X"20203135"; -- 015
							 l <= 3;
			 when X"10" =>  A <= X"20203136"; -- 016
							 l <= 3;
			 when X"11" =>  A <= X"20203137"; -- 017
							 l <= 3;
			 when X"12" =>  A <= X"20203138"; -- 018
							 l <= 3;
			 when X"13" =>  A <= X"20203139"; -- 019
							 l <= 3;
			 when X"14" =>  A <= X"20203230"; -- 020
							 l <= 3;
			 when X"15" =>  A <= X"20203231"; -- 021
							 l <= 3;
			 when X"16" =>  A <= X"20203232"; -- 022
							 l <= 3;
			 when X"17" =>  A <= X"20203233"; -- 023
							 l <= 3;
			 when X"18" =>  A <= X"20203234"; -- 024
							 l <= 3;
			 when X"19" =>  A <= X"20203235"; -- 025
							 l <= 3;
			 when X"1a" =>  A <= X"20203236"; -- 026
							 l <= 3;
			 when X"1b" =>  A <= X"20203237"; -- 027
							 l <= 3;
			 when X"1c" =>  A <= X"20203238"; -- 028
							 l <= 3;
			 when X"1d" =>  A <= X"20203239"; -- 029
							 l <= 3;
			 when X"1e" =>  A <= X"20203330"; -- 030
							 l <= 3;
			 when X"1f" =>  A <= X"20203331"; -- 031
							 l <= 3;
			 when X"20" =>  A <= X"20203332"; -- 032
							 l <= 3;
			 when X"21" =>  A <= X"20203333"; -- 033
							 l <= 3;
			 when X"22" =>  A <= X"20203334"; -- 034
							 l <= 3;
			 when X"23" =>  A <= X"20203335"; -- 035
							 l <= 3;
			 when X"24" =>  A <= X"20203336"; -- 036
							 l <= 3;
			 when X"25" =>  A <= X"20203337"; -- 037
							 l <= 3;
			 when X"26" =>  A <= X"20203338"; -- 038
							 l <= 3;
			 when X"27" =>  A <= X"20203339"; -- 039
							 l <= 3;
			 when X"28" =>  A <= X"20203430"; -- 040
							 l <= 3;
			 when X"29" =>  A <= X"20203431"; -- 041
							 l <= 3;
			 when X"2a" =>  A <= X"20203432"; -- 042
							 l <= 3;
			 when X"2b" =>  A <= X"20203433"; -- 043
							 l <= 3;
			 when X"2c" =>  A <= X"20203434"; -- 044
							 l <= 3;
			 when X"2d" =>  A <= X"20203435"; -- 045
							 l <= 3;
			 when X"2e" =>  A <= X"20203436"; -- 046
							 l <= 3;
			 when X"2f" =>  A <= X"20203437"; -- 047
							 l <= 3;
			 when X"30" =>  A <= X"20203438"; -- 048
							 l <= 3;
			 when X"31" =>  A <= X"20203439"; -- 049
							 l <= 3;
			 when X"32" =>  A <= X"20203530"; -- 050
							 l <= 3;
			 when X"33" =>  A <= X"20203531"; -- 051
							 l <= 3;
			 when X"34" =>  A <= X"20203532"; -- 052
							 l <= 3;
			 when X"35" =>  A <= X"20203533"; -- 053
							 l <= 3;
			 when X"36" =>  A <= X"20203534"; -- 054
							 l <= 3;
			 when X"37" =>  A <= X"20203535"; -- 055
							 l <= 3;
			 when X"38" =>  A <= X"20203536"; -- 056
							 l <= 3;
			 when X"39" =>  A <= X"20203537"; -- 057
							 l <= 3;
			 when X"3a" =>  A <= X"20203538"; -- 058
							 l <= 3;
			 when X"3b" =>  A <= X"20203539"; -- 059
							 l <= 3;
			 when X"3c" =>  A <= X"20203630"; -- 060
							 l <= 3;
			 when X"3d" =>  A <= X"20203631"; -- 061
							 l <= 3;
			 when X"3e" =>  A <= X"20203632"; -- 062
							 l <= 3;
			 when X"3f" =>  A <= X"20203633"; -- 063
							 l <= 3;
			 when X"40" =>  A <= X"20203634"; -- 064
							 l <= 3;
			 when X"41" =>  A <= X"20203635"; -- 065
							 l <= 3;
			 when X"42" =>  A <= X"20203636"; -- 066
							 l <= 3;
			 when X"43" =>  A <= X"20203637"; -- 067
							 l <= 3;
			 when X"44" =>  A <= X"20203638"; -- 068
							 l <= 3;
			 when X"45" =>  A <= X"20203639"; -- 069
							 l <= 3;
			 when X"46" =>  A <= X"20203730"; -- 070
							 l <= 3;
			 when X"47" =>  A <= X"20203731"; -- 071
							 l <= 3;
			 when X"48" =>  A <= X"20203732"; -- 072
							 l <= 3;
			 when X"49" =>  A <= X"20203733"; -- 073
							 l <= 3;
			 when X"4a" =>  A <= X"20203734"; -- 074
							 l <= 3;
			 when X"4b" =>  A <= X"20203735"; -- 075
							 l <= 3;
			 when X"4c" =>  A <= X"20203736"; -- 076
							 l <= 3;
			 when X"4d" =>  A <= X"20203737"; -- 077
							 l <= 3;
			 when X"4e" =>  A <= X"20203738"; -- 078
							 l <= 3;
			 when X"4f" =>  A <= X"20203739"; -- 079
							 l <= 3;
			 when X"50" =>  A <= X"20203830"; -- 080
							 l <= 3;
			 when X"51" =>  A <= X"20203831"; -- 081
							 l <= 3;
			 when X"52" =>  A <= X"20203832"; -- 082
							 l <= 3;
			 when X"53" =>  A <= X"20203833"; -- 083
							 l <= 3;
			 when X"54" =>  A <= X"20203834"; -- 084
							 l <= 3;
			 when X"55" =>  A <= X"20203835"; -- 085
							 l <= 3;
			 when X"56" =>  A <= X"20203836"; -- 086
							 l <= 3;
			 when X"57" =>  A <= X"20203837"; -- 087
							 l <= 3;
			 when X"58" =>  A <= X"20203838"; -- 088
							 l <= 3;
			 when X"59" =>  A <= X"20203839"; -- 089
							 l <= 3;
			 when X"5a" =>  A <= X"20203930"; -- 090
							 l <= 3;
			 when X"5b" =>  A <= X"20203931"; -- 091
							 l <= 3;
			 when X"5c" =>  A <= X"20203932"; -- 092
							 l <= 3;
			 when X"5d" =>  A <= X"20203933"; -- 093
							 l <= 3;
			 when X"5e" =>  A <= X"20203934"; -- 094
							 l <= 3;
			 when X"5f" =>  A <= X"20203935"; -- 095
							 l <= 3;
			 when X"60" =>  A <= X"20203936"; -- 096
							 l <= 3;
			 when X"61" =>  A <= X"20203937"; -- 097
							 l <= 3;
			 when X"62" =>  A <= X"20203938"; -- 098
							 l <= 3;
			 when X"63" =>  A <= X"20203939"; -- 099
							 l <= 3;
			 when X"64" =>  A <= X"20313030"; -- 100
							 l <= 4;
			 when X"65" =>  A <= X"20313031"; -- 101
							 l <= 4;
			 when X"66" =>  A <= X"20313032"; -- 102
							 l <= 4;
			 when X"67" =>  A <= X"20313033"; -- 103
							 l <= 4;
			 when X"68" =>  A <= X"20313034"; -- 104
							 l <= 4;
			 when X"69" =>  A <= X"20313035"; -- 105
							 l <= 4;
			 when X"6a" =>  A <= X"20313036"; -- 106
							 l <= 4;
			 when X"6b" =>  A <= X"20313037"; -- 107
							 l <= 4;
			 when X"6c" =>  A <= X"20313038"; -- 108
							 l <= 4;
			 when X"6d" =>  A <= X"20313039"; -- 109
							 l <= 4;
			 when X"6e" =>  A <= X"20313130"; -- 110
							 l <= 4;
			 when X"6f" =>  A <= X"20313131"; -- 111
							 l <= 4;
			 when X"70" =>  A <= X"20313132"; -- 112
							 l <= 4;
			 when X"71" =>  A <= X"20313133"; -- 113
							 l <= 4;
			 when X"72" =>  A <= X"20313134"; -- 114
							 l <= 4;
			 when X"73" =>  A <= X"20313135"; -- 115
							 l <= 4;
			 when X"74" =>  A <= X"20313136"; -- 116
							 l <= 4;
			 when X"75" =>  A <= X"20313137"; -- 117
							 l <= 4;
			 when X"76" =>  A <= X"20313138"; -- 118
							 l <= 4;
			 when X"77" =>  A <= X"20313139"; -- 119
							 l <= 4;
			 when X"78" =>  A <= X"20313230"; -- 120
							 l <= 4;
			 when X"79" =>  A <= X"20313231"; -- 121
							 l <= 4;
			 when X"7a" =>  A <= X"20313232"; -- 122
							 l <= 4;
			 when X"7b" =>  A <= X"20313233"; -- 123
							 l <= 4;
			 when X"7c" =>  A <= X"20313234"; -- 124
							 l <= 4;
			 when X"7d" =>  A <= X"20313235"; -- 125
							 l <= 4;
			 when X"7e" =>  A <= X"20313236"; -- 126
							 l <= 4;
			 when X"7f" =>  A <= X"20313237"; -- 127
							 l <= 4;
			 when X"80" =>  A <= X"20313238"; -- 128
							 l <= 4;
			 when X"81" =>  A <= X"20313239"; -- 129
							 l <= 4;
			 when X"82" =>  A <= X"20313330"; -- 130
							 l <= 4;
			 when X"83" =>  A <= X"20313331"; -- 131
							 l <= 4;
			 when X"84" =>  A <= X"20313332"; -- 132
							 l <= 4;
			 when X"85" =>  A <= X"20313333"; -- 133
							 l <= 4;
			 when X"86" =>  A <= X"20313334"; -- 134
							 l <= 4;
			 when X"87" =>  A <= X"20313335"; -- 135
							 l <= 4;
			 when X"88" =>  A <= X"20313336"; -- 136
							 l <= 4;
			 when X"89" =>  A <= X"20313337"; -- 137
							 l <= 4;
			 when X"8a" =>  A <= X"20313338"; -- 138
							 l <= 4;
			 when X"8b" =>  A <= X"20313339"; -- 139
							 l <= 4;
			 when X"8c" =>  A <= X"20313430"; -- 140
							 l <= 4;
			 when X"8d" =>  A <= X"20313431"; -- 141
							 l <= 4;
			 when X"8e" =>  A <= X"20313432"; -- 142
							 l <= 4;
			 when X"8f" =>  A <= X"20313433"; -- 143
							 l <= 4;
			 when X"90" =>  A <= X"20313434"; -- 144
							 l <= 4;
			 when X"91" =>  A <= X"20313435"; -- 145
							 l <= 4;
			 when X"92" =>  A <= X"20313436"; -- 146
							 l <= 4;
			 when X"93" =>  A <= X"20313437"; -- 147
							 l <= 4;
			 when X"94" =>  A <= X"20313438"; -- 148
							 l <= 4;
			 when X"95" =>  A <= X"20313439"; -- 149
							 l <= 4;
			 when X"96" =>  A <= X"20313530"; -- 150
							 l <= 4;
			 when X"97" =>  A <= X"20313531"; -- 151
							 l <= 4;
			 when X"98" =>  A <= X"20313532"; -- 152
							 l <= 4;
			 when X"99" =>  A <= X"20313533"; -- 153
							 l <= 4;
			 when X"9a" =>  A <= X"20313534"; -- 154
							 l <= 4;
			 when X"9b" =>  A <= X"20313535"; -- 155
							 l <= 4;
			 when X"9c" =>  A <= X"20313536"; -- 156
							 l <= 4;
			 when X"9d" =>  A <= X"20313537"; -- 157
							 l <= 4;
			 when X"9e" =>  A <= X"20313538"; -- 158
							 l <= 4;
			 when X"9f" =>  A <= X"20313539"; -- 159
							 l <= 4;
			 when X"a0" =>  A <= X"20313630"; -- 160
							 l <= 4;
			 when X"a1" =>  A <= X"20313631"; -- 161
							 l <= 4;
			 when X"a2" =>  A <= X"20313632"; -- 162
							 l <= 4;
			 when X"a3" =>  A <= X"20313633"; -- 163
							 l <= 4;
			 when X"a4" =>  A <= X"20313634"; -- 164
							 l <= 4;
			 when X"a5" =>  A <= X"20313635"; -- 165
							 l <= 4;
			 when X"a6" =>  A <= X"20313636"; -- 166
							 l <= 4;
			 when X"a7" =>  A <= X"20313637"; -- 167
							 l <= 4;
			 when X"a8" =>  A <= X"20313638"; -- 168
							 l <= 4;
			 when X"a9" =>  A <= X"20313639"; -- 169
							 l <= 4;
			 when X"aa" =>  A <= X"20313730"; -- 170
							 l <= 4;
			 when X"ab" =>  A <= X"20313731"; -- 171
							 l <= 4;
			 when X"ac" =>  A <= X"20313732"; -- 172
							 l <= 4;
			 when X"ad" =>  A <= X"20313733"; -- 173
							 l <= 4;
			 when X"ae" =>  A <= X"20313734"; -- 174
							 l <= 4;
			 when X"af" =>  A <= X"20313735"; -- 175
							 l <= 4;
			 when X"b0" =>  A <= X"20313736"; -- 176
							 l <= 4;
			 when X"b1" =>  A <= X"20313737"; -- 177
							 l <= 4;
			 when X"b2" =>  A <= X"20313738"; -- 178
							 l <= 4;
			 when X"b3" =>  A <= X"20313739"; -- 179
							 l <= 4;
			 when X"b4" =>  A <= X"20313830"; -- 180
							 l <= 4;
			 when X"b5" =>  A <= X"20313831"; -- 181
							 l <= 4;
			 when X"b6" =>  A <= X"20313832"; -- 182
							 l <= 4;
			 when X"b7" =>  A <= X"20313833"; -- 183
							 l <= 4;
			 when X"b8" =>  A <= X"20313834"; -- 184
							 l <= 4;
			 when X"b9" =>  A <= X"20313835"; -- 185
							 l <= 4;
			 when X"ba" =>  A <= X"20313836"; -- 186
							 l <= 4;
			 when X"bb" =>  A <= X"20313837"; -- 187
							 l <= 4;
			 when X"bc" =>  A <= X"20313838"; -- 188
							 l <= 4;
			 when X"bd" =>  A <= X"20313839"; -- 189
							 l <= 4;
			 when X"be" =>  A <= X"20313930"; -- 190
							 l <= 4;
			 when X"bf" =>  A <= X"20313931"; -- 191
							 l <= 4;
			 when X"c0" =>  A <= X"20313932"; -- 192
							 l <= 4;
			 when X"c1" =>  A <= X"20313933"; -- 193
							 l <= 4;
			 when X"c2" =>  A <= X"20313934"; -- 194
							 l <= 4;
			 when X"c3" =>  A <= X"20313935"; -- 195
							 l <= 4;
			 when X"c4" =>  A <= X"20313936"; -- 196
							 l <= 4;
			 when X"c5" =>  A <= X"20313937"; -- 197
							 l <= 4;
			 when X"c6" =>  A <= X"20313938"; -- 198
							 l <= 4;
			 when X"c7" =>  A <= X"20313939"; -- 199
							 l <= 4;
			 when X"c8" =>  A <= X"20323030"; -- 200
							 l <= 4;
			 when X"c9" =>  A <= X"20323031"; -- 201
							 l <= 4;
			 when X"ca" =>  A <= X"20323032"; -- 202
							 l <= 4;
			 when X"cb" =>  A <= X"20323033"; -- 203
							 l <= 4;
			 when X"cc" =>  A <= X"20323034"; -- 204
							 l <= 4;
			 when X"cd" =>  A <= X"20323035"; -- 205
							 l <= 4;
			 when X"ce" =>  A <= X"20323036"; -- 206
							 l <= 4;
			 when X"cf" =>  A <= X"20323037"; -- 207
							 l <= 4;
			 when X"d0" =>  A <= X"20323038"; -- 208
							 l <= 4;
			 when X"d1" =>  A <= X"20323039"; -- 209
							 l <= 4;
			 when X"d2" =>  A <= X"20323130"; -- 210
							 l <= 4;
			 when X"d3" =>  A <= X"20323131"; -- 211
							 l <= 4;
			 when X"d4" =>  A <= X"20323132"; -- 212
							 l <= 4;
			 when X"d5" =>  A <= X"20323133"; -- 213
							 l <= 4;
			 when X"d6" =>  A <= X"20323134"; -- 214
							 l <= 4;
			 when X"d7" =>  A <= X"20323135"; -- 215
							 l <= 4;
			 when X"d8" =>  A <= X"20323136"; -- 216
							 l <= 4;
			 when X"d9" =>  A <= X"20323137"; -- 217
							 l <= 4;
			 when X"da" =>  A <= X"20323138"; -- 218
							 l <= 4;
			 when X"db" =>  A <= X"20323139"; -- 219
							 l <= 4;
			 when X"dc" =>  A <= X"20323230"; -- 220
							 l <= 4;
			 when X"dd" =>  A <= X"20323231"; -- 221
							 l <= 4;
			 when X"de" =>  A <= X"20323232"; -- 222
							 l <= 4;
			 when X"df" =>  A <= X"20323233"; -- 223
							 l <= 4;
			 when X"e0" =>  A <= X"20323234"; -- 224
							 l <= 4;
			 when X"e1" =>  A <= X"20323235"; -- 225
							 l <= 4;
			 when X"e2" =>  A <= X"20323236"; -- 226
							 l <= 4;
			 when X"e3" =>  A <= X"20323237"; -- 227
							 l <= 4;
			 when X"e4" =>  A <= X"20323238"; -- 228
							 l <= 4;
			 when X"e5" =>  A <= X"20323239"; -- 229
							 l <= 4;
			 when X"e6" =>  A <= X"20323330"; -- 230
							 l <= 4;
			 when X"e7" =>  A <= X"20323331"; -- 231
							 l <= 4;
			 when X"e8" =>  A <= X"20323332"; -- 232
							 l <= 4;
			 when X"e9" =>  A <= X"20323333"; -- 233
							 l <= 4;
			 when X"ea" =>  A <= X"20323334"; -- 234
							 l <= 4;
			 when X"eb" =>  A <= X"20323335"; -- 235
							 l <= 4;
			 when X"ec" =>  A <= X"20323336"; -- 236
							 l <= 4;
			 when X"ed" =>  A <= X"20323337"; -- 237
							 l <= 4;
			 when X"ee" =>  A <= X"20323338"; -- 238
							 l <= 4;
			 when X"ef" =>  A <= X"20323339"; -- 239
							 l <= 4;
			 when X"f0" =>  A <= X"20323430"; -- 240
							 l <= 4;
			 when X"f1" =>  A <= X"20323431"; -- 241
							 l <= 4;
			 when X"f2" =>  A <= X"20323432"; -- 242
							 l <= 4;
			 when X"f3" =>  A <= X"20323433"; -- 243
							 l <= 4;
			 when X"f4" =>  A <= X"20323434"; -- 244
							 l <= 4;
			 when X"f5" =>  A <= X"20323435"; -- 245
							 l <= 4;
			 when X"f6" =>  A <= X"20323436"; -- 246
							 l <= 4;
			 when X"f7" =>  A <= X"20323437"; -- 247
							 l <= 4;
			 when X"f8" =>  A <= X"20323438"; -- 248
							 l <= 4;
			 when X"f9" =>  A <= X"20323439"; -- 249
							 l <= 4;
			 when X"fa" =>  A <= X"20323530"; -- 250
							 l <= 4;
			 when X"fb" =>  A <= X"20323531"; -- 251
							 l <= 4;
			 when X"fc" =>  A <= X"20323532"; -- 252
							 l <= 4;
			 when X"fd" =>  A <= X"20323533"; -- 253
							 l <= 4;
			 when X"fe" =>  A <= X"20323534"; -- 254
							 l <= 4;
			 when X"ff" =>  A <= X"20323535"; -- 255
							 l <= 4;
			 when others => 
		end case;
end process;


end Behavioral;

